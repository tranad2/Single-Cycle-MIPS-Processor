LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY pipeMW IS
	PORT (
		clk: IN STD_LOGIC;
		WB_in: IN STD_LOGIC;
		WriteRegM: IN STD_LOGIC;
		ReadDataM: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		ALUInM: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		WB_out: OUT STD_LOGIC;
		WriteRegW: IN STD_LOGIC;
		ReadDataW: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		ALUOutW: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END pipeMW;

ARCHITECTURE arch_pipe of pipeMW IS
BEGIN

END arch_pipe;