LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY pipeFD IS
	PORT (
		clk: IN STD_LOGIC;
		FlushE: IN STD_LOGIC;
		rdata_1_in: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		rdata_2_in: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		RsD: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		RtD: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		RdD: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		SignImmD: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		rdata_1_out: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		rdata_2_out: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		RsE: OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		RtE: OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		RdE: OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		SignImmE: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	);
END pipeFD;

ARCHITECTURE arch_pipe of pipeFD IS
BEGIN

END arch_pipe;