LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY pipeFD IS
	PORT (
		clk: IN STD_LOGIC;
		stallF: IN STD_LOGIC;
		PC_in: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		PC_out: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END pipeFD;

ARCHITECTURE arch_pipe of pipeFD IS
BEGIN

END arch_pipe;